package FirstAttempt;
String s = "Hello World";
module mkAttempt;
endmodule
endpackage