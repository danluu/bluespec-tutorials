package FirstAttempt;
String s = "Hello World";
endpackage