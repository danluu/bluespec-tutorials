package TL0;

interface TL;
endinterface: TL

module sysTL(TL);
endmodule: sysTL

endpackage: TL0

