package FirstAttempt;
	//huzzah!
endpackage